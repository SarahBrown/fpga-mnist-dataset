module sevenSeg(
	input[3:0] sel,
	output[7:0]segs);
	
	assign segs = 	(sel == 4'h0) ? 8'b11000000:
						(sel == 4'h1) ? 8'b11111001:
						(sel == 4'h2) ? 8'b10100100:
						(sel == 4'h3) ? 8'b10110000:
						(sel == 4'h4) ? 8'b10011001:
						(sel == 4'h5) ? 8'b10010010:
						(sel == 4'h6) ? 8'b10000010:
						(sel == 4'h7) ? 8'b11111000:
						(sel == 4'h8) ? 8'b10000000:
						(sel == 4'h9) ? 8'b10011000:
						(sel == 4'ha) ? 8'b10001000:
						(sel == 4'hb) ? 8'b10000011:
						(sel == 4'hc) ? 8'b11000110:
						(sel == 4'hd) ? 8'b10100001:
						(sel == 4'he) ? 8'b10000110:
						(sel == 4'hf) ? 8'b00001110:
											 8'b11111111;
endmodule